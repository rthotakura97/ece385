module font_rom ( input [7:0]	addr,
		  output [7:0]	data
					 );

	parameter ADDR_WIDTH = 8;
   	parameter DATA_WIDTH =  8;
	logic [ADDR_WIDTH-1:0] addr_reg;
				
	// ROM definition				
	parameter [0:2**ADDR_WIDTH-1][DATA_WIDTH-1:0] ROM = {

         // code x00
        8'b00000000, // 0
        8'b00000000, // 1
        8'b01111100, // 2  *****
        8'b11000110, // 3 **   **
        8'b11000110, // 4 **   **
        8'b11001110, // 5 **  ***
        8'b11011110, // 6 ** ****
        8'b11110110, // 7 **** **
        8'b11100110, // 8 ***  **
        8'b11000110, // 9 **   **
        8'b11000110, // a **   **
        8'b01111100, // b  *****
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x01
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00011000, // 2
        8'b00111000, // 3
        8'b01111000, // 4    **
        8'b00011000, // 5   ***
        8'b00011000, // 6  ****
        8'b00011000, // 7    **
        8'b00011000, // 8    **
        8'b00011000, // 9    **
        8'b00011000, // a    **
        8'b01111110, // b    **
        8'b00000000, // c    **
        8'b00000000, // d  ******
        8'b00000000, // e
        8'b00000000, // f
         // code x02
        8'b00000000, // 0
        8'b00000000, // 1
        8'b01111100, // 2  *****
        8'b11000110, // 3 **   **
        8'b00000110, // 4      **
        8'b00001100, // 5     **
        8'b00011000, // 6    **
        8'b00110000, // 7   **
        8'b01100000, // 8  **
        8'b11000000, // 9 **
        8'b11000110, // a **   **
        8'b11111110, // b *******
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x03
        8'b00000000, // 0
        8'b00000000, // 1
        8'b01111100, // 2  *****
        8'b11000110, // 3 **   **
        8'b00000110, // 4      **
        8'b00000110, // 5      **
        8'b00111100, // 6   ****
        8'b00000110, // 7      **
        8'b00000110, // 8      **
        8'b00000110, // 9      **
        8'b11000110, // a **   **
        8'b01111100, // b  *****
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x04
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00001100, // 2     **
        8'b00011100, // 3    ***
        8'b00111100, // 4   ****
        8'b01101100, // 5  ** **
        8'b11001100, // 6 **  **
        8'b11111110, // 7 *******
        8'b00001100, // 8     **
        8'b00001100, // 9     **
        8'b00001100, // a     **
        8'b00011110, // b    ****
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x05
        8'b00000000, // 0
        8'b00000000, // 1
        8'b11111110, // 2 *******
        8'b11000000, // 3 **
        8'b11000000, // 4 **
        8'b11000000, // 5 **
        8'b11111100, // 6 ******
        8'b00000110, // 7      **
        8'b00000110, // 8      **
        8'b00000110, // 9      **
        8'b11000110, // a **   **
        8'b01111100, // b  *****
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x06
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00111000, // 2   ***
        8'b01100000, // 3  **
        8'b11000000, // 4 **
        8'b11000000, // 5 **
        8'b11111100, // 6 ******
        8'b11000110, // 7 **   **
        8'b11000110, // 8 **   **
        8'b11000110, // 9 **   **
        8'b11000110, // a **   **
        8'b01111100, // b  *****
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x07
        8'b00000000, // 0
        8'b00000000, // 1
        8'b11111110, // 2 *******
        8'b11000110, // 3 **   **
        8'b00000110, // 4      **
        8'b00000110, // 5      **
        8'b00001100, // 6     **
        8'b00011000, // 7    **
        8'b00110000, // 8   **
        8'b00110000, // 9   **
        8'b00110000, // a   **
        8'b00110000, // b   **
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x08
        8'b00000000, // 0
        8'b00000000, // 1
        8'b01111100, // 2  *****
        8'b11000110, // 3 **   **
        8'b11000110, // 4 **   **
        8'b11000110, // 5 **   **
        8'b01111100, // 6  *****
        8'b11000110, // 7 **   **
        8'b11000110, // 8 **   **
        8'b11000110, // 9 **   **
        8'b11000110, // a **   **
        8'b01111100, // b  *****
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x09
        8'b00000000, // 0
        8'b00000000, // 1
        8'b01111100, // 2  *****
        8'b11000110, // 3 **   **
        8'b11000110, // 4 **   **
        8'b11000110, // 5 **   **
        8'b01111110, // 6  ******
        8'b00000110, // 7      **
        8'b00000110, // 8      **
        8'b00000110, // 9      **
        8'b00001100, // a     **
        8'b01111000, // b  ****
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
        // Unused
        8'b00000000,
        8'b00000000,
        8'b00000000, 
        8'b00000000, 
        8'b00000000, 
        8'b00000000, 
        8'b00000000, 
        8'b00000000, 
        8'b00000000, 
        8'b00000000, 
        8'b00000000, 
        8'b00000000, 
        8'b00000000, 
        8'b00000000, 
        8'b00000000, 
        8'b00000000,
 
        8'b00000000,
        8'b00000000,
        8'b00000000, 
        8'b00000000, 
        8'b00000000, 
        8'b00000000, 
        8'b00000000, 
        8'b00000000, 
        8'b00000000, 
        8'b00000000, 
        8'b00000000, 
        8'b00000000, 
        8'b00000000, 
        8'b00000000, 
        8'b00000000, 
        8'b00000000,
 
        8'b00000000,
        8'b00000000,
        8'b00000000, 
        8'b00000000, 
        8'b00000000, 
        8'b00000000, 
        8'b00000000, 
        8'b00000000, 
        8'b00000000, 
        8'b00000000, 
        8'b00000000, 
        8'b00000000, 
        8'b00000000, 
        8'b00000000, 
        8'b00000000, 
        8'b00000000,
 
        8'b00000000,
        8'b00000000,
        8'b00000000, 
        8'b00000000, 
        8'b00000000, 
        8'b00000000, 
        8'b00000000, 
        8'b00000000, 
        8'b00000000, 
        8'b00000000, 
        8'b00000000, 
        8'b00000000, 
        8'b00000000, 
        8'b00000000, 
        8'b00000000, 
        8'b00000000,
 
        8'b00000000,
        8'b00000000,
        8'b00000000, 
        8'b00000000, 
        8'b00000000, 
        8'b00000000, 
        8'b00000000, 
        8'b00000000, 
        8'b00000000, 
        8'b00000000, 
        8'b00000000, 
        8'b00000000, 
        8'b00000000, 
        8'b00000000, 
        8'b00000000, 
        8'b00000000, 
        8'b00000000,

        8'b00000000,
        8'b00000000, 
        8'b00000000, 
        8'b00000000, 
        8'b00000000, 
        8'b00000000, 
        8'b00000000, 
        8'b00000000, 
        8'b00000000, 
        8'b00000000, 
        8'b00000000, 
        8'b00000000, 
        8'b00000000, 
        8'b00000000, 
        8'b00000000, 
        };

	assign data = ROM[addr];

endmodule  
